LIBRARY ieee ;
 USE ieee.std_logic_1164.all ;
ENTITY DECOMOD IS
 PORT ( w : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		en:IN STD_LOGIC; 
 y : OUT STD_LOGIC_VECTOR(15 DOWNTO 0) ) ; 
 END DECOMOD ;
ARCHITECTURE Behavior OF DECOMOD IS 
 signal x : STD_LOGIC_VECTOR(2 DOWNTO 0) ; 
 BEGIN x <= en & w;
  WITH x SELECT 
 
 y <= "0000000000000001" WHEN "0000",
 "0000000000000010" WHEN "0001",
 "0000000000000100" WHEN "0010",
 "0000000000001000" WHEN "0011",
 "0000000000010000" WHEN "0100",
 "0000000000100000" WHEN "0101",
 "0000000001000000" WHEN "0110",
 "0000000010000000" WHEN "0111",
 
 
 "0000000100000000" WHEN "1000",
 "0000001000000000" WHEN "1001",
 "0000010000000000" WHEN "1010",
 "0000100000000000" WHEN "1011",
 "0001000000000000" WHEN "1100",
 "0010000000000000" WHEN "1101",
 "0100000000000000" WHEN "1110",
 "1000000000000000" WHEN "1111";

 

 END Behavior ;